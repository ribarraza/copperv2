interface copperv2_bfm;
    bit         bus_ir_addr_ready;
    wire        bus_ir_addr_valid;
    wire [31:0] bus_ir_addr_bits;
    wire        bus_ir_data_ready;
    bit         bus_ir_data_valid;
    bit  [31:0] bus_ir_data_bits;
    bit         bus_dr_addr_ready;
    wire        bus_dr_addr_valid;
    wire [31:0] bus_dr_addr_bits;
    wire        bus_dr_data_ready;
    bit         bus_dr_data_valid;
    bit  [31:0] bus_dr_data_bits;
    bit         bus_dw_req_ready;
    wire        bus_dw_req_valid;
    wire [31:0] bus_dw_req_bits_data;
    wire [31:0] bus_dw_req_bits_addr;
    wire [7:0]  bus_dw_req_bits_strobe;
    wire        bus_dw_resp_ready;
    bit         bus_dw_resp_valid;
    bit         bus_dw_resp_bits;

//   assign op = op_set;
//
//   task reset_alu();
//      reset_n = 1'b0;
//      @(negedge clk);
//      @(negedge clk);
//      reset_n = 1'b1;
//      start = 1'b0;
//   endtask : reset_alu
//   
//
//
//   task send_op(input byte iA, input byte iB, input operation_t iop, output shortint alu_result);
//      if (iop == rst_op) begin
//         @(posedge clk);
//         reset_n = 1'b0;
//         start = 1'b0;
//         @(posedge clk);
//         #1;
//         reset_n = 1'b1;
//      end else begin
//         @(negedge clk);
//         op_set = iop;
//         A = iA;
//         B = iB;
//         start = 1'b1;
//         if (iop == no_op) begin
//            @(posedge clk);
//            #1;
//            start = 1'b0;           
//         end else begin
//            do
//              @(negedge clk);
//            while (done == 0);
//            alu_result = result;
//            start = 1'b0;
//         end
//      end // else: !if(iop == rst_op)
//      
//   endtask : send_op
//   
//   command_monitor command_monitor_h;
//
//   function operation_t op2enum();
//      case(op)
//        3'b000 : return no_op;
//        3'b001 : return add_op;
//        3'b010 : return and_op;
//        3'b011 : return xor_op;
//        3'b100 : return mul_op;
//        default : $fatal("Illegal operation on op bus");
//      endcase // case (op)
//   endfunction : op2enum
//
//
//   always @(posedge clk) begin : op_monitor
//      static bit in_command = 0;
//      if (start) begin : start_high
//        if (!in_command) begin : new_command
//           command_monitor_h.write_to_monitor(A, B, op2enum());
//           in_command = (op2enum() != no_op);
//        end : new_command
//      end : start_high
//      else // start low
//        in_command = 0;
//   end : op_monitor
//
//   always @(negedge reset_n) begin : rst_monitor
//      if (command_monitor_h != null) //guard against VCS time 0 negedge
//        command_monitor_h.write_to_monitor($random,0,rst_op);
//   end : rst_monitor
//   
//   result_monitor  result_monitor_h;
//
//   initial begin : result_monitor_thread
//      forever begin : result_monitor_block
//         @(posedge clk) ;
//         if (done) 
//           result_monitor_h.write_to_monitor(result);
//      end : result_monitor_block
//   end : result_monitor_thread
//   
//
//   initial begin
//      clk = 0;
//      fork
//         forever begin
//            #10;
//            clk = ~clk;
//         end
//      join_none
//   end
//

endinterface : copperv2_bfm
